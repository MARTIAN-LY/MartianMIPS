`include "define.vh"


module martianmips (
    input   wire    clk,
    input   wire    rst
);

endmodule //martianmips