`include "define.vh"


module martianmips (
    input   wire    clk,
    input   wire    rst,

    input   wire[`RegBus]
);

endmodule //martianmips