`include "define.vh"



module regfile (
    input   wire    clk,
    input   wire    rst,

    //写端口
    input   wire    we,                 //写使能
    input   wire[`RegAddBus]    waddr,  //写地址
    input   wire[`RegBus]


);

endmodule //regfile