module id (
    input   wire    rst,
    
);

endmodule //id